
module cpulyc (
	probe,
	source);	

	input	[0:0]	probe;
	output	[0:0]	source;
endmodule
